// AlarmClockHDL_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module AlarmClockHDL_tb (
	);

	wire        alarmclockhdl_inst_clk_bfm_clk_clk;            // AlarmClockHDL_inst_clk_bfm:clk -> AlarmClockHDL_inst:clk_clk
	wire  [0:0] alarmclockhdl_inst_alarm1_bfm_conduit_export;  // AlarmClockHDL_inst_alarm1_bfm:sig_export -> AlarmClockHDL_inst:alarm1_export
	wire  [0:0] alarmclockhdl_inst_button1_bfm_conduit_export; // AlarmClockHDL_inst_button1_bfm:sig_export -> AlarmClockHDL_inst:button1_export
	wire  [0:0] alarmclockhdl_inst_button2_bfm_conduit_export; // AlarmClockHDL_inst_button2_bfm:sig_export -> AlarmClockHDL_inst:button2_export
	wire  [0:0] alarmclockhdl_inst_button3_bfm_conduit_export; // AlarmClockHDL_inst_button3_bfm:sig_export -> AlarmClockHDL_inst:button3_export
	wire  [0:0] alarmclockhdl_inst_button4_bfm_conduit_export; // AlarmClockHDL_inst_button4_bfm:sig_export -> AlarmClockHDL_inst:button4_export
	wire  [1:0] alarmclockhdl_inst_buzzer_export;              // AlarmClockHDL_inst:buzzer_export -> AlarmClockHDL_inst_buzzer_bfm:sig_export
	wire  [6:0] alarmclockhdl_inst_segment1_export;            // AlarmClockHDL_inst:segment1_export -> AlarmClockHDL_inst_segment1_bfm:sig_export
	wire  [6:0] alarmclockhdl_inst_segment2_export;            // AlarmClockHDL_inst:segment2_export -> AlarmClockHDL_inst_segment2_bfm:sig_export
	wire  [6:0] alarmclockhdl_inst_segment3_export;            // AlarmClockHDL_inst:segment3_export -> AlarmClockHDL_inst_segment3_bfm:sig_export
	wire  [6:0] alarmclockhdl_inst_segment4_export;            // AlarmClockHDL_inst:segment4_export -> AlarmClockHDL_inst_segment4_bfm:sig_export

	AlarmClockHDL alarmclockhdl_inst (
		.alarm1_export   (alarmclockhdl_inst_alarm1_bfm_conduit_export),  //   alarm1.export
		.button1_export  (alarmclockhdl_inst_button1_bfm_conduit_export), //  button1.export
		.button2_export  (alarmclockhdl_inst_button2_bfm_conduit_export), //  button2.export
		.button3_export  (alarmclockhdl_inst_button3_bfm_conduit_export), //  button3.export
		.button4_export  (alarmclockhdl_inst_button4_bfm_conduit_export), //  button4.export
		.buzzer_export   (alarmclockhdl_inst_buzzer_export),              //   buzzer.export
		.clk_clk         (alarmclockhdl_inst_clk_bfm_clk_clk),            //      clk.clk
		.segment1_export (alarmclockhdl_inst_segment1_export),            // segment1.export
		.segment2_export (alarmclockhdl_inst_segment2_export),            // segment2.export
		.segment3_export (alarmclockhdl_inst_segment3_export),            // segment3.export
		.segment4_export (alarmclockhdl_inst_segment4_export)             // segment4.export
	);

	altera_conduit_bfm alarmclockhdl_inst_alarm1_bfm (
		.sig_export (alarmclockhdl_inst_alarm1_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm alarmclockhdl_inst_button1_bfm (
		.sig_export (alarmclockhdl_inst_button1_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm alarmclockhdl_inst_button2_bfm (
		.sig_export (alarmclockhdl_inst_button2_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm alarmclockhdl_inst_button3_bfm (
		.sig_export (alarmclockhdl_inst_button3_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm alarmclockhdl_inst_button4_bfm (
		.sig_export (alarmclockhdl_inst_button4_bfm_conduit_export)  // conduit.export
	);

	altera_conduit_bfm_0002 alarmclockhdl_inst_buzzer_bfm (
		.sig_export (alarmclockhdl_inst_buzzer_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) alarmclockhdl_inst_clk_bfm (
		.clk (alarmclockhdl_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0003 alarmclockhdl_inst_segment1_bfm (
		.sig_export (alarmclockhdl_inst_segment1_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarmclockhdl_inst_segment2_bfm (
		.sig_export (alarmclockhdl_inst_segment2_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarmclockhdl_inst_segment3_bfm (
		.sig_export (alarmclockhdl_inst_segment3_export)  // conduit.export
	);

	altera_conduit_bfm_0003 alarmclockhdl_inst_segment4_bfm (
		.sig_export (alarmclockhdl_inst_segment4_export)  // conduit.export
	);

endmodule
